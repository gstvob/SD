library ieee;
use ieee.std_logic_1164.all;

entity decod7seg is
port( inpt : in std_logic_vector(3 downto 0);
		outp : out std_logic_vector(6 downto 0)
);
end;

architecture decod7seg_behv of decod7seg is
begin

--decodificador basico que simplesmente pega uma entrada de 4 bits e transforma para um display de 7 segmentos.
	with inpt select
		outp <= "1111001" when "0001",
				  "0100100" when "0010",
				  "0110000" when "0011",
				  "0011001" when "0100",
				  "0010010" when "0101",
				  "0000010" when "0110",
				  "1111000" when "0111",
				  "0000000" when "1000",
				  "0010000" when "1001",
				  "1000000" when others;
end;
